package shared_pkg;
    logic test_finished;
    int error_cnt, correct_cnt;
    event emonitor;
endpackage
